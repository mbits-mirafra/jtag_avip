`ifndef JTAGCONTROLLERDEVICEPATTERNBASEDVIRTUALSEQUENCE_INCLUDED_
`define JTAGCONTROLLERDEVICEPATTERNBASEDVIRTUALSEQUENCE_INCLUDED_

class JtagVirtualControllerDevicePatternBasedSequence extends JtagVirtualBaseSequence;
  `uvm_object_utils(JtagVirtualControllerDevicePatternBasedSequence)

  JtagControllerDevicePatternBasedSequence jtagControllerDevicePatternBasedSequence;
  JtagTargetDeviceBaseSequence  jtagTargetDeviceBaseSequence;
  JtagControllerDeviceAgentConfig jtagControllerDeviceAgentConfig;

  extern function new(string name = "JtagVirtualControllerDevicePatternBasedSequence");
  extern virtual task body();
  extern task setConfig(JtagControllerDeviceAgentConfig jtagControllerDeviceAgentConfig);
endclass : JtagVirtualControllerDevicePatternBasedSequence 


function JtagControllerDevicePatternBasedVirtualSequence ::new(string name = "JtagVirtualControllerDevicePatternBasedSequence");
  super.new(name);
endfunction  : new

task JtagControllerDevicePatternBasedVirtualSequence :: body();
  super.body();
  `uvm_do_on_with(jtagControllerDevicePatternBasedSequence,p_sequencer.jtagControllerDeviceSequencer,{patternNeeded == jtagControllerDeviceAgentConfig.patternNeeded;})
endtask : body 

task JtagControllerDevicePatternBasedVirtualSequence :: setConfig(JtagControllerDeviceAgentConfig jtagControllerDeviceAgentConfig);
  this.jtagControllerDeviceAgentConfig = jtagControllerDeviceAgentConfig;
endtask : setConfig
 
`endif
