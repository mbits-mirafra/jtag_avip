`ifndef JTAGTDIWidth32INSTRUCTIONWIDTH4TEST_INCLUDED_
`define JTAGTDIWidth32INSTRUCTIONWIDTH4TEST_INCLUDED_

class JtagTdiWidth32InstructionWidth4Test extends JtagBaseTest;
  `uvm_component_utils( JtagTdiWidth32InstructionWidth4Test)

  extern function new(string name = "JtagTdiWidth32InstructionWidth4Test" , uvm_component parent);
  extern virtual function void build_phase(uvm_phase phase);
  extern virtual task run_phase (uvm_phase phase);
endclass :  JtagTdiWidth32InstructionWidth4Test

function  JtagTdiWidth32InstructionWidth4Test :: new(string name = "JtagTdiWidth32InstructionWidth4Test" , uvm_component parent);
  super.new(name,parent);
endfunction : new

function void JtagTdiWidth32InstructionWidth4Test :: build_phase(uvm_phase phase);
  super.build_phase(phase);
  jtagEnvConfig.jtagControllerDeviceAgentConfig.jtagTestVectorWidth = testVectorWidth32Bit;
  jtagEnvConfig.jtagControllerDeviceAgentConfig.jtagInstructionWidth = instructionWidth4Bit;
  jtagEnvConfig.jtagTargetDeviceAgentConfig.jtagTestVectorWidth = testVectorWidth32Bit;
  jtagEnvConfig.jtagTargetDeviceAgentConfig.jtagInstructionWidth = instructionWidth4Bit;
endfunction : build_phase

task JtagTdiWidth32InstructionWidth4Test :: run_phase(uvm_phase phase);
  jtagVirtualControllerDeviceTestingSequence = JtagVirtualControllerDeviceTestingSequence :: type_id :: create("jtagVirtualControllerDeviceTestingSequence");
  jtagVirtualControllerDeviceTestingSequence.setConfig(jtagEnvConfig.jtagControllerDeviceAgentConfig);
 
  phase.raise_objection(this);
  repeat( NO_OF_TESTS) begin 
    jtagVirtualControllerDeviceTestingSequence.start(jtagEnv.jtagVirtualSequencer);
  end 
  phase.drop_objection(this);

endtask : run_phase

`endif
